module turnOnLED (output led);

/* Turn-on LED */ 
assign led = 1'b0;

endmodule
